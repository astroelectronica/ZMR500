.title KiCad schematic
.include "C:/AE/ZMR500/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/ZMR500/_models/C3216X5R1C106M160AA_p.mod"
.include "C:/AE/ZMR500/_models/C3216X7R2A105M160AA_p.mod"
.include "C:/AE/ZMR500/_models/ZMR500.spice.txt"
XU5 /VOUT 0 C2012X7R2A104K125AA_p
XU3 /VIN 0 C2012X7R2A104K125AA_p
I1 /VOUT 0 {ILOAD}
V1 /VIN 0 {VSOURCE}
XU1 /VIN 0 /VOUT ZMR500
XU2 /VIN 0 C3216X7R2A105M160AA_p
XU4 /VOUT 0 C3216X5R1C106M160AA_p
.end
